`timescale 1 ns / 1 ps
module READ_ROM32 ( input[4:0] ADDR ,output[31:0] DATA_RE,output[31:0] DATA_IM);
reg [31:0] re[0:31];
initial  begin
re[0] = 32'h00000000;re[1] = 32'hFFE4CC88;re[2] = 32'h002DA5B3;re[3] = 32'hFFCE9932;
re[4] = 32'h00254173;re[5] = 32'hFFF2E19A;re[6] = 32'hFFF0C26D;re[7] = 32'h0026B1CD;
re[8] = 32'hFFCE4E3A;re[9] = 32'h002CB328;re[10] = 32'hFFE6AE85;re[11] = 32'hFFFDC9B2;
re[12] = 32'h001D07D3;re[13] = 32'hFFD17EA5;re[14] = 32'h00310311;re[15] = 32'hFFDC4195;
re[16] = 32'h000AF8A5;re[17] = 32'h0011551D;re[18] = 32'hFFD7F13F;re[19] = 32'h0031E3D5;
re[20] = 32'hFFD455CB;re[21] = 32'h001762CC;re[22] = 32'h00046B81;re[23] = 32'hFFE13261;
re[24] = 32'h002F45B3;re[25] = 32'hFFCF793E;re[26] = 32'h00222978;re[27] = 32'hFFF7329D;
re[28] = 32'hFFEC9C0A;re[29] = 32'h002957A0;re[30] = 32'hFFCE0320;re[31] = 32'h002A8B5D;
end
reg [31:0] im[0:31];
initial  begin
im[0] = 32'h00000000;im[1] = 32'h00000000;im[2] = 32'h00000000;im[3] = 32'h00000000;
im[4] = 32'h00000000;im[5] = 32'h00000000;im[6] = 32'h00000000;im[7] = 32'h00000000;
im[8] = 32'h00000000;im[9] = 32'h00000000;im[10] = 32'h00000000;im[11] = 32'h00000000;
im[12] = 32'h00000000;im[13] = 32'h00000000;im[14] = 32'h00000000;im[15] = 32'h00000000;
im[16] = 32'h00000000;im[17] = 32'h00000000;im[18] = 32'h00000000;im[19] = 32'h00000000;
im[20] = 32'h00000000;im[21] = 32'h00000000;im[22] = 32'h00000000;im[23] = 32'h00000000;
im[24] = 32'h00000000;im[25] = 32'h00000000;im[26] = 32'h00000000;im[27] = 32'h00000000;
im[28] = 32'h00000000;im[29] = 32'h00000000;im[30] = 32'h00000000;im[31] = 32'h00000000;
end
assign DATA_RE = re[ADDR];
assign DATA_IM = im[ADDR];
endmodule